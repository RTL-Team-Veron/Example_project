package rtl_pkg;
	parameter DW = 4;
endpackage
